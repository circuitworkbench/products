.TITLE cccs
V1 1 GND 20.0
R1 1 2 2.4
R2 3 GND 1.333
//CCCS F1
VF1 2 3
F1 GND 3 VF1 200m
.OP
.END